`include "../00_bench/agent/and_agent/and_if.sv"  
`include "../00_bench/agent/and_agent/and_agent.sv"
