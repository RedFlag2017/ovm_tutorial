`include "../03_testcase/tc01/tc01.sv"