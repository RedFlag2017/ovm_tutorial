`include "../00_bench/testbench/tb.sv"